library verilog;
use verilog.vl_types.all;
entity brainfuck_cpu_tb is
end brainfuck_cpu_tb;
